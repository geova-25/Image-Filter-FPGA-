module InstructionMemory2(
    input wire  [31:0] DIR,
    output reg [31:0] DO
    );
	 
	
	 always@(*)
	 begin
			case (DIR)
				32'h00000000: DO <= 32'h0F000000;
				32'h00000004: DO <= 32'h0F000000;
				32'h00000008: DO <= 32'h0F000000;
				32'h0000000C: DO <= 32'h0F000000;
				32'h00000010: DO <= 32'hED000000;
				32'h00000014: DO <= 32'h0F000000;
				32'h00000018: DO <= 32'h0F000000;
				32'h0000001C: DO <= 32'hED100004;
				32'h00000020: DO <=32'h7D200028;
				32'h00000024: DO <=32'h7D300001;
				32'h00000028: DO <=32'h7D400000;
				32'h0000002C: DO <=32'h4C510000;
				32'h00000030: DO <=32'h1D640005;
				32'h00000034: DO <=32'h4C730000;
				32'h00000038: DO <=32'h8C065000;
				32'h0000003C: DO <=32'h92000013;
				32'h00000040: DO <=32'h0F000000;
				32'h00000044: DO <=32'h0F000000;
				32'h00000048: DO <=32'h0CB42000;
				32'h0000004C: DO <=32'hAC0B0000;
				32'h00000050: DO <=32'h0F000000;
				32'h00000054: DO <=32'h0F000000;
				32'h00000058: DO <=32'hBC900000;
				32'h0000005C: DO <=32'h1DAB0002;
				32'h00000060: DO <=32'h0F000000;
				32'h00000064: DO <=32'h0F000000;
				32'h00000068: DO <=32'hFC0A9000;
				32'h0000006C: DO <=32'h8C067000;
				32'h00000070: DO <=32'h15440004;
				32'h00000074: DO <=32'h15330001;
				32'h00000078: DO <=32'h0F000000;
				32'h0000007C: DO <=32'h0F000000;
				32'h00000080: DO <=32'h19440001;
				32'h00000084: DO <=32'h9EFFFFE9;
				32'h00000088: DO <=32'h0F000000;
				32'h0000008C: DO <=32'h0F000000;
				32'h00000090: DO <=32'h9EFFFFFE;
				32'h00000094: DO <=32'h0F000000;
				32'h00000098: DO <=32'h0F000000;
				default:  	  DO <=32'h0F000000;
			endcase
	 end

 /*
always@(*)
	 begin
			case (DIR)
				32'h00000000: DO <= 32'h0F000000;
				32'h00000004: DO <= 32'h0F000000;
				32'h00000008: DO <= 32'h0F000000;
				32'h0000000C: DO <= 32'h0F000000;
				32'h00000010: DO <= 32'hED000000;
				32'h00000014: DO <= 32'h0F000000;
				32'h00000018: DO <= 32'h0F000000;
				32'h0000001C: DO <= 32'hED100004;
				32'h00000020: DO <=32'h7D200028;
				32'h00000024: DO <=32'h7D300001;
				32'h00000028: DO <=32'h7D400000;
				32'h0000002C: DO <=32'h4C510000;
				32'h00000030: DO <=32'h1D640005;
				32'h00000034: DO <=32'h4C730000;
				32'h00000038: DO <=32'h8C065000;
				32'h0000003C: DO <=32'h92000013;
				32'h00000040: DO <=32'h0F000000;
				32'h00000044: DO <=32'h0F000000;
				32'h00000048: DO <=32'h0CB42000;
				32'h0000004C: DO <=32'hAC0B0000;
				32'h00000050: DO <=32'h0F000000;
				32'h00000054: DO <=32'h0F000000;
				32'h00000058: DO <=32'hBC900000;
				32'h0000005C: DO <=32'h1DAB0002;
				32'h00000060: DO <=32'h0F000000;
				32'h00000064: DO <=32'h0F000000;
				32'h00000068: DO <=32'hFC0A9000;
				32'h0000006C: DO <=32'h8C067000;
				32'h00000070: DO <=32'h15440004;
				32'h00000074: DO <=32'h15330001;
				32'h00000078: DO <=32'h0F000000;
				32'h0000007C: DO <=32'h0F000000;
				32'h00000080: DO <=32'h19440001;
				32'h00000084: DO <=32'h9EFFFFE9;
				32'h00000088: DO <=32'h0F000000;
				32'h0000008C: DO <=32'h0F000000;
				
				32'h00000090: DO <=32'h7D400000;
				32'h00000094: DO <=32'h8C040000;
				32'h00000098: DO <=32'h0F000000;
				32'h0000009C: DO <=32'h0F000000;
				32'h000000A0: DO <=32'h9600003A;
				32'h000000A4: DO <=32'h7D300000;
				32'h000000A8: DO <=32'h3D610002;
				32'h000000AC: DO <=32'h8C036000;
				32'h000000B0: DO <=32'h0F000000;
				32'h000000B4: DO <=32'h0F000000;
				32'h000000B8: DO <=32'h96000030;
				32'h000000BC: DO <=32'h0C742000;
				32'h000000C0: DO <=32'h4C830000;
				32'h000000C4: DO <=32'h3D880003;
				32'h000000C8: DO <=32'h0C887000;
				32'h000000CC: DO <=32'hCC880000;
				32'h000000D0: DO <=32'hED900008;
				32'h000000D4: DO <=32'h0F000000;
				32'h000000D8: DO <=32'h5C889000;
				32'h000000DC: DO <=32'h1D930001;
				32'h000000E0: DO <=32'h4C990000;
				32'h000000E4: DO <=32'h3D990002;
				32'h000000E8: DO <=32'h0C979000;
				32'h000000EC: DO <=32'h0F000000;
				32'h000000F0: DO <=32'hCC990000;
				32'h000000F4: DO <=32'hEDA0000C;
				32'h000000F8: DO <=32'h0F000000;
				32'h000000FC: DO <=32'h5C99A000;
				32'h00000100: DO <=32'h1DA30002;
				32'h00000104: DO <=32'h4CA0A000;
				32'h00000108: DO <=32'h3DAA0001;
				32'h0000010C: DO <=32'h0CDA7000;
				32'h00000110: DO <=32'hCCAD0000;
				32'h00000114: DO <=32'hEDB0000A;
				32'h00000118: DO <=32'h0F000000;
				32'h0000011C: DO <=32'h5CAAB000;
				32'h00000120: DO <=32'h1DB30003;
				32'h00000124: DO <=32'h4CBB0000;
				32'h00000128: DO <=32'h0CBB7000;
				32'h0000012C: DO <=32'hCCBB0000;
				32'h00000130: DO <=32'hEDC00014;
				32'h00000134: DO <=32'h0F000000;
				32'h00000138: DO <=32'h5CBBC000;
				32'h0000013C: DO <=32'h1DF30004;
				32'h00000140: DO <=32'h4CFF0000;
				32'h00000144: DO <=32'h0CFF7000;
				32'h00000148: DO <=32'hCCFF0000;
				32'h0000014C: DO <=32'h0F000000;
				32'h00000150: DO <=32'h5CFF0000;
				32'h00000154: DO <=32'h6CE89000;
				32'h00000158: DO <=32'h6CEEA000;
				32'h0000015C: DO <=32'h6CEEB000;
				32'h00000160: DO <=32'h1D330001;
				32'h00000164: DO <=32'hBC800000;
				32'h00000168: DO <=32'h0F000000;
				32'h0000016C: DO <=32'h0F000000;
				32'h00000170: DO <=32'hFC0D8000;
				32'h00000174: DO <=32'h0F000000;
				32'h00000178: DO <=32'h0F000000;
				32'h0000017C: DO <=32'h9EFFFFC9;
				32'h00000180: DO <=32'h1D440001;
				32'h00000184: DO <=32'h0F000000;
				32'h00000188: DO <=32'h0F000000;
				32'h0000018C: DO <=32'h9EFFFFC0;
				32'h00000190: DO <=32'h0F000000;
				32'h00000194: DO <=32'h0F000000;
				32'h00000198: DO <=32'h9EFFFFE6;
				32'h0000019C: DO <= 32'h0F000000;
				32'h00000200: DO <= 32'h0F000000;
								
				
				
				default:  	  DO <=32'h0F000000;
			endcase
			
	 end*/


	 
endmodule