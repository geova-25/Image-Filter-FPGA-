module InstructionMemory2(
    input wire  [31:0] DIR,
    output reg [31:0] DO
    );
	 
	 
	 always@(*)
	 begin
			case (DIR)
				32'h00000000: DO <= 32'h0F000000;
				32'h00000004: DO <= 32'h0F000000;
				32'h00000008: DO <= 32'h0F000000;
				32'h0000000C: DO <= 32'h0F000000;
				32'h00000010: DO <= 32'hED000000;
				32'h00000014: DO <= 32'h0F000000;
				32'h00000018: DO <= 32'h0F000000;
				32'h0000001C: DO <= 32'hED100004;
				32'h00000020: DO <=32'h7D200028;
				32'h00000024: DO <=32'h7D300001;
				32'h00000028: DO <=32'h7D400000;
				32'h0000002C: DO <=32'h4C510000;
				32'h00000030: DO <=32'h1D640005;
				32'h00000034: DO <=32'h4C730000;
				32'h00000038: DO <=32'h8C065000;
				32'h0000003C: DO <=32'h92000013;
				32'h00000040: DO <=32'h0F000000;
				32'h00000044: DO <=32'h0F000000;
				32'h00000048: DO <=32'h0CB42000;
				32'h0000004C: DO <=32'hAC0B0000;
				32'h00000050: DO <=32'h0F000000;
				32'h00000054: DO <=32'h0F000000;
				32'h00000058: DO <=32'hBC900000;
				32'h0000005C: DO <=32'h1DAB0002;
				32'h00000060: DO <=32'h0F000000;
				32'h00000064: DO <=32'h0F000000;
				32'h00000068: DO <=32'hFC0A9000;
				32'h0000006C: DO <=32'h8C067000;
				32'h00000070: DO <=32'h15440004;
				32'h00000074: DO <=32'h15330001;
				32'h00000078: DO <=32'h0F000000;
				32'h0000007C: DO <=32'h0F000000;
				32'h00000080: DO <=32'h19440001;
				32'h00000084: DO <=32'h9EFFFFE9;
				32'h00000088: DO <=32'h0F000000;
				32'h0000008C: DO <=32'h0F000000;
				32'h00000090: DO <=32'h9EFFFFFE;
				32'h00000094: DO <=32'h0F000000;
				32'h00000098: DO <=32'h0F000000;
				default:  	  DO <=32'h0F000000;
			endcase
	 end


	 
endmodule